LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY DRAKES_DATA_PATH IS
GENERIC( P:INTEGER:=64;
	 MW:INTEGER:=128;
	 E: INTEGER:= 128;
	 M: INTEGER:= 128
);

-- GLOBAL CONTROL VALUES

PORT(
	CLK: IN STD_LOGIC;
	RESET: IN STD_LOGIC;
	PRODUCT_REG_EN: IN STD_LOGIC;
	ALU_SEL: IN STD_LOGIC_VECTOR(1 downto 0);
	MCAND_REG_EN: IN STD_LOGIC;
	MULT_REG_EN: IN STD_LOGIC

);
END DRAKES_DATA_PATH;


ARCHITECTURE STRUCTURAL OF DRAKES_DATA_PATH is



-- ALU --
COMPONENT DRAKES_ALU is 
generic( width: natural := 64;
	output: natural	:= 128);
port(
	alu_in1: in std_logic_vector(output-1 downto 0);
	alu_in2: in std_logic_vector(output-1 downto 0);
	alu_sel: in std_logic_vector(1 downto 0);
	alu_out: out std_logic_vector(output-1 downto 0)
);
end COMPONENT;


-- MCAND LEFT SHIFT REGISTER

COMPONENT shift_LEFT_128BIT is 
generic( width: NATURAL);
port(	
		CLK: IN STD_LOGIC;
		RST: IN STD_LOGIC;
		EN: IN STD_LOGIC;
		OP_Q: out std_logic_vector(width-1 downto 0)
	);
end COMPONENT;


-- MULT SHIFT RIGHT VALUES

COMPONENT shift_RIGHT_64BIT is 
generic( width: NATURAL);
port(	
		CLK: IN STD_LOGIC;
		RST: IN STD_LOGIC;
		EN: IN STD_LOGIC;
		OP_Q: out std_logic_vector(width-1 downto 0)
	);
end COMPONENT;


-- PRODUCT REGISTER 

COMPONENT Drakes_PRODUCT_Reg is

	GENERIC(
		P :integer:= 128);	
	 PORT(	
		CLK: IN STD_LOGIC;
		RST: IN STD_LOGIC;
		EN: IN STD_LOGIC;
		OP_A: IN STD_LOGIC_VECTOR(P-1 DOWNTO 0);
		OP_Q: OUT STD_LOGIC_VECTOR(P-1 DOWNTO 0));
	END COMPONENT;



----------------------------------
-- 			SIGNALS				--
----------------------------------


SIGNAL ALU_OUT: STD_LOGIC_VECTOR(MW-1 DOWNTO 0);
SIGNAL PRODUCT_REG_OUT: STD_LOGIC_VECTOR(MW-1 DOWNTO 0);
SIGNAL MCAND_REG_OUT: STD_LOGIC_VECTOR(MW-1 DOWNTO 0);
SIGNAL MULT_REG_OUT: STD_LOGIC_VECTOR(P-1 DOWNTO 0);

BEGIN

I1_ALU: DRAKES_ALU GENERIC MAP(P,MW)PORT MAP(PRODUCT_REG_OUT, MCAND_REG_OUT, ALU_SEL, ALU_OUT);
I2_PRODUCT_REG: DRAKES_PRODUCT_REG GENERIC MAP(MW)PORT MAP(CLK, RESET, MULT_REG_OUT(0), ALU_OUT, PRODUCT_REG_OUT);
I3_MCAND_REG: shift_LEFT_128BIT GENERIC MAP(MW)PORT MAP(CLK, RESET, MCAND_REG_EN, MCAND_REG_OUT);
I4_MULT_REG: shift_RIGHT_64BIT GENERIC MAP(P)PORT MAP(CLK, RESET, MULT_REG_EN,  MULT_REG_OUT);


END STRUCTURAL;