LIBRARY IEEE;
USE work.CLOCKS.all;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_textio.all;
USE std.textio.all;
USE work.txt_util.all;

ENTITY tb_MULTIPLIER IS
END;

ARCHITECTURE TESTBENCH OF tb_MULTIPLIER is

CONSTANT P: INTEGER:=64;
CONSTANT MW: INTEGER:=128;



COMPONENT DRAKES_MULTIPLIER_DATAPATH

GENERIC(    P: INTEGER:=64;
            MW: INTEGER:=128);

PORT(

    CLK: IN STD_LOGIC;
	RESET: IN STD_LOGIC;
	PRODUCT_REG_EN: IN STD_LOGIC;
	ALU_SEL: IN STD_LOGIC_VECTOR(1 downto 0);
	MCAND_REG_EN: IN STD_LOGIC;
	MULT_REG_EN: IN STD_LOGIC;
	MULT_DIRECTION: IN STD_LOGIC;
	MCAND_DIRECTION: IN STD_LOGIC
    
);

END COMPONENT;



BEGIN



END TESTBENCH;